library verilog;
use verilog.vl_types.all;
entity CPU_TB is
end CPU_TB;
