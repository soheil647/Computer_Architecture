library verilog;
use verilog.vl_types.all;
entity CPU_TEST is
end CPU_TEST;
