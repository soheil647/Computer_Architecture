library verilog;
use verilog.vl_types.all;
entity Stack_tb is
end Stack_tb;
