library verilog;
use verilog.vl_types.all;
entity exp_controller is
    generic(
        \IF\            : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        \TOS\           : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        JUMP            : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        JUMPZ           : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        PUSH1           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        PUSH2           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        POP1            : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        POP2            : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        POP3            : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        Rtype0          : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1);
        Rtype1          : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi0);
        Rtype2          : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1);
        RtypeNOT        : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi0);
        RtypeEND        : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi1);
        ADD             : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        SUB             : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        \AND\           : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        \NOT\           : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        \PUSH\          : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        \POP\           : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        JMP             : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        JZ              : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1)
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        Opcode          : in     vl_logic_vector(2 downto 0);
        IorD            : out    vl_logic;
        MtoS            : out    vl_logic;
        srcA            : out    vl_logic;
        srcB            : out    vl_logic;
        PCwrite         : out    vl_logic;
        PCwritecond     : out    vl_logic;
        PCsrc           : out    vl_logic;
        IRwrite         : out    vl_logic;
        MemRead         : out    vl_logic;
        MemWrite        : out    vl_logic;
        ldA             : out    vl_logic;
        ldB             : out    vl_logic;
        push            : out    vl_logic;
        pop             : out    vl_logic;
        tos             : out    vl_logic;
        ALUOperation    : out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of \IF\ : constant is 1;
    attribute mti_svvh_generic_type of \TOS\ : constant is 1;
    attribute mti_svvh_generic_type of JUMP : constant is 1;
    attribute mti_svvh_generic_type of JUMPZ : constant is 1;
    attribute mti_svvh_generic_type of PUSH1 : constant is 1;
    attribute mti_svvh_generic_type of PUSH2 : constant is 1;
    attribute mti_svvh_generic_type of POP1 : constant is 1;
    attribute mti_svvh_generic_type of POP2 : constant is 1;
    attribute mti_svvh_generic_type of POP3 : constant is 1;
    attribute mti_svvh_generic_type of Rtype0 : constant is 1;
    attribute mti_svvh_generic_type of Rtype1 : constant is 1;
    attribute mti_svvh_generic_type of Rtype2 : constant is 1;
    attribute mti_svvh_generic_type of RtypeNOT : constant is 1;
    attribute mti_svvh_generic_type of RtypeEND : constant is 1;
    attribute mti_svvh_generic_type of ADD : constant is 1;
    attribute mti_svvh_generic_type of SUB : constant is 1;
    attribute mti_svvh_generic_type of \AND\ : constant is 1;
    attribute mti_svvh_generic_type of \NOT\ : constant is 1;
    attribute mti_svvh_generic_type of \PUSH\ : constant is 1;
    attribute mti_svvh_generic_type of \POP\ : constant is 1;
    attribute mti_svvh_generic_type of JMP : constant is 1;
    attribute mti_svvh_generic_type of JZ : constant is 1;
end exp_controller;
